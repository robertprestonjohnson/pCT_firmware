//Complete DAQ program for six chips, to run in the FPGA on the pCTFE64 test board.
//To be increased to 12 chips when a complete board is available.
//This version leaves the trigger decisions to the event builder FPGA.
//R. Johnson     Rewrite in March 2013 to simplify commands that had evolved over time.
//Modified June 10, 2013 to remove the buffer clear signal.  Added local check for buffer overwrite.

module FPGA_DAQ_TKR6(Dout,FastOR,CMDtoChips,Tack,Clock,ResetHard,CmdIn,TrgIn,Data,TReq,Address);
input [3:0] Address;  //FPGA address, on the tracker boards to be set by dip switches
input Clock;          //Clock for the FPGA (C9, A9)    (Phase-shifted output clock needs to go to P8, T8 to send clock to the chips)
input ResetHard;      //Reset everything, including the command decoding state machine (P7, M7)
input CmdIn;          //Input DAQ commands (F7, E6)
input TrgIn;          //Tack input (D5, C5)
input [5:0] Data;     //Serial data streams from the pCTFE64 chips (B15, B16) (F12, G11) (D14, D16) (F13, F14) (C15, C16) (E15, E16)
input [5:0] TReq;     //Trigger outputs from the pCTFE64 chips (M5, N4) (R2, R1) (P2, P1) (N3, N1) (M2, M1) (L3, L1)
output Tack;          //Trigger acknowledge going to the pCTFE64 chips (M9, N8)
output CMDtoChips;    //Commands going to the pCTFE64 chips (R9, T9)
output Dout;          //Output serial data stream (B6, A6)
output FastOR;        //Output OR of all 6 trigger requests (B5, A5)

wire [5:0] Data,TReq;
wire [3:0] Address;
reg Dout, CMDtoChips;

reg CalStrobe;			//Signal that a calibration command has been sent to the ASICs
reg Reset;    			//Reset pulse generated by command
wire [3:0] UnDoBuf;    	//Signal that the corresponding front-end buffer has cleared

reg Parity;			//Parity calculated for local command received 
reg Error;			//Store parity error
reg [9:0] CmdSav;   //Saved ASIC command string, extracted from the incoming bit stream
reg InProg;			//Set while a run is in progress
reg EndRun;			//Pulse to signal end of run
reg [5:0] StrtSq;   //Start sequence for register readback, inserted before the bits from the ASIC

reg MuxData, SendEvt;
reg [77:0] RegOut;	//Register for shifting out the test string and DAQ counters

//Command definitions (3-bit commands to this FPGA program)
// 0: Send a test string back to the DAQ
// 1: Unused
// 2: Start a run.  During the run, no commands should be sent except for read and end-run.  
// 3: End a run.
// 4: Read back parity error bit and DAQ counters
//    This will also clear the parity error flag, unless this command generates a new error.
// 5: Reset counters and variables in this code
// 6: Reset the front-end ASICs without altering their registers (takes about 1 millisecond to complete)
// 7: Read a merged event from the local buffers and send it to the event builder (as soon as it is available)

//Command format:
//  start bit
//  4-bit address of the FPGA board
//  routing bit:  1=complete command to ASICs follows    0=command to this program
//  3-bit local command  
//  parity bit, not counting the start bit
//
//	Note:  during a run no commands should be sent besides end-run (except that Read commands will be
//         sent automatically from the event builder buffer manager).  This program is not protected against
//         receiving other commands, such as read register, which would disrupt the data acquisition.  To avoid
//         delaying the data acquisition, the incoming commands stream is not checked before forwarding it to 
//         the ASICs.  This program also does not check the parity of ASIC commands.  But the ASICs themselves
//         will do that.

initial begin
//	$display("Time     StateTOT TReqChip CalStrobe CntStrt CntTOT CntShft TOTHeader TOTNclus MuxData");
//  $display("Time        State    CmdIn TrgIn   Cnt   InProg Data   TReq CMD Dout RegIn   StrtSq TC RRC StateRd CntRd2 TrgCode RdStrng SndEvt");
end

always @ (posedge Clock) begin
//   $display("%g\t  %b %b     %b  %b %b   %b %b %b   %b       %b %b %b %b %b     %b    %b  %b    %b",$time,State,CmdIn,TrgIn, Cnt,InProg,Data,TReq,CMDtoChips,Dout,RegIn,StrtSq,ThisFPGA,ReadRegCmd,StateRd,CntRd2,TrgCode,RdString,SendEvt);
end

assign Tack = TrgIn;   //Pass the trigger acknowledge straight through to the ASICs
assign TReqChip =   TReq[0] | TReq[1] | TReq[2] | TReq[3] | TReq[4] | TReq[5];
assign FastOR =  InProg & TReqChip;  //Tracker self triggering
always @ (posedge FastOR) $display("%g\t FPGA_DAQ %d:  FastOR fires;  TReq=%b",$time,Address,TReq);

//Count triggers
reg [31:0] Ntriggers;
reg [15:0] NReads, NSends;
wire [1:0] TrgTag;
reg [3:0] BufOcc;
reg TrgErr;
TriggerReceiver_RTL TrigDecode(Clock,ResetHard,TrgIn,TrgPls,TrgTag);
always @ (posedge Clock) begin
	if (Reset) begin
		Ntriggers <= 0;
		BufOcc <= 4'b0000;
		TrgErr <= 1'b0;
	end else begin
		if (TrgPls) begin
			Ntriggers <= Ntriggers + 1;
			if (!UnDoBuf[TrgTag]) BufOcc[TrgTag] <= 1'b1;
			if (BufOcc[TrgTag]) TrgErr <= 1'b1;
		end else begin
			if (UnDoBuf[TrgTag]) BufOcc[TrgTag] <= 1'b0;
		end
	end
end

//Names given to the eight commands:
parameter cmdTest = 3'b000;
parameter cmdFeCd = 3'b001;
parameter cmdStRn = 3'b010;
parameter cmdEnRn = 3'b011;
parameter cmdRdFg = 3'b100;
parameter cmdRset = 3'b101;
parameter cmdRsCh = 3'b110;
parameter cmdSend = 3'b111;

//State machine to interpret and execute commands sent from the event builder
//Encoding of states:
parameter [10:0] Wait = 11'b00000000001;  //Wait for a start bit
parameter [10:0] RdBt = 11'b00000000010;  //Read the 4-bit address
parameter [10:0] Brch = 11'b00000000100;  //Branch to chip vs local command
parameter [10:0] ACmd = 11'b00000001000;  //Clock in the ASIC command and start bit
parameter [10:0] FeCd = 11'b00000010000;  //Check the ASIC command
parameter [10:0] Ct66 = 11'b00000100000;  //Wait some more clock cycles for the command to end or register data to come back
parameter [10:0] RdCm = 11'b00001000000;  //Read in the 3-bit local command
parameter [10:0] Deco = 11'b00010000000;  //Decode the local command
parameter [10:0] Prty = 11'b00100000000;  //Check parity of local command
parameter [10:0] WrWd = 11'b01000000000;  //Write out monitoring information or a test string
parameter [10:0] WtDn = 11'b10000000000;  //Wait for front-end reset to finish

reg [10:0] State, NextState;
reg [7:0] Cnt;     	//Eight-bit counter
reg [2:0] RegIn;   	//Register for shifting in and storing the command 
reg [3:0] AddrIn;   //Register for shifting in the FPGA address
reg [6:0] nDat;   	//Number of clocks needed to complete a front-end ASIC command
reg ResetSlow;

always @ (State or CmdIn or Cnt or DoneRst or InProg or nDat or RegIn)
begin:CombinatorialLogic
  case(State)
	Wait: 	begin
				if (CmdIn == 1'b1)   	//Trigger state machine on command start bit
					NextState=RdBt;
				else
					NextState=Wait;
			end
	RdBt:	begin
				if (Cnt == 3)			//Count in four address bits
					NextState=Brch;
				else
					NextState=RdBt;
			end
	Brch:	begin						//Branch to ASIC command or local command
				if (CmdIn) NextState=ACmd;
				else NextState=RdCm;
			end
	ACmd:	begin
			    if (Cnt == 9)			//Count in five ASIC address bits and 4 command bits
					NextState=FeCd;
				else
					NextState=ACmd;
			end
	FeCd:	begin
				NextState=Ct66;			//Look at the command received and set nDat; direct bit stream to ASICs
			end
	Ct66:	begin
				if (Cnt[6:0] == nDat)	//Wait long enough for command bits to go to ASIC and register data to come back
					NextState=Wait;
				else
					NextState=Ct66;
			end
	RdCm:	begin
				if (Cnt == 2) NextState = Deco;		//Count in the 3 local command bits
				else NextState = RdCm;
			end
	Deco:   begin
				case (RegIn)						//Branch to appropriate execution for the command received
					cmdTest: NextState = WrWd;
					cmdFeCd: NextState = Prty;   //Do nothing
					cmdStRn: NextState = Prty;
					cmdEnRn: NextState = Prty;
					cmdRdFg: if (InProg)
								NextState=Prty;
							 else
								NextState=WrWd;
					cmdRset: NextState = Prty;
					cmdRsCh: NextState = WtDn;  
					cmdSend: NextState = Prty;
				endcase
			end
	WtDn:	begin								//Wait for the complete reset of the ASICs to complete (about 1 millisecond)
				if (DoneRst) NextState=Prty;
				else NextState=WtDn;
			end
	Prty:	begin								//Check the parity of the received local command (should be positive)
				NextState=Wait;
			end
	WrWd:	begin								//Shift a test string or DAQ counters into the output data stream
				if (Cnt==77)
					NextState=Prty;
				else
					NextState=WrWd;
			end
	default:begin
				NextState=Wait;
			end
  endcase
 end
 
always @ (posedge Clock)
begin:SequentialLogic
  if (Reset) begin				//This Reset is activated by command, but also by the ResetHard
	Error <= 1'b0;
	NReads <= 0;
	NSends <= 0;
	SendEvt <= 1'b0;
	InProg <= 1'b0;
	EndRun <= 1'b0;
	CalStrobe <= 1'b0;
  end
  if (ResetHard) begin			//This reset is received from the event builder over a dedicated link
	Reset <= 1'b1;
	ResetSlow <= 1'b0;
	State <= Wait;
  end else begin
    State <= NextState;
	case(State)
		Wait: 	begin
					Reset <= 1'b0;
					Cnt <= 0;
					Parity <= 1'b0; 
				end
		RdBt:	begin
					Cnt <= Cnt + 1;
					Parity <= Parity^CmdIn;     	//Calculate parity of the incoming address and command bits
					AddrIn <= {AddrIn[2:0],CmdIn};	//Shift in the 4-bit FPGA address of the incoming command
				end
		Brch:	begin
//					$display("%g\t FPGA_DAQ %d:  received command for address %b, branch to %b",$time,Address,AddrIn,CmdIn);
					Cnt <= 0;
				end
		ACmd:	begin
//					$display("%g\t FPGA_DAQ %d:  %b CMDtoChips=%b,  Dout=%b",$time,Address,State,CMDtoChips,Dout);
					Cnt <= Cnt + 1;
					CmdSav <= {CmdSav[8:0],CmdIn};	//Shift in the 5-bit ASIC address and 4-bit command
				end
		FeCd:	begin
//					$display("%g\t FPGA_DAQ_TKR6:  %b CMDtoChips=%b,  Dout=%b",$time,State,CMDtoChips,Dout);
//					$display("%g\t FPGA_DAQ %d:  ASIC command code = %b, Chip %d, Command=%h",$time,Address,CmdSav,CmdSav[8:4],CmdSav[3:0]);
					Cnt <= 0;
					case (CmdSav[3:0])      //Set the length of the data field or returned data as appropriate for each command
						4'h0: nDat <= 0;
						4'h1: begin nDat <= 0; $display("%g\t FPGA_DAQ_TKR6: soft reset going to chips.",$time); end
						4'h2: begin nDat <= 1; NReads <= NReads + 1; end  
						4'h3: begin nDat <= 71;  StrtSq <= {2'b11,Address}; end
						4'h4: begin nDat <= 71;  StrtSq <= {2'b11,Address}; end
						4'h5: begin nDat <= 71;  StrtSq <= {2'b11,Address}; end
						4'h6: begin nDat <= 71;  StrtSq <= {2'b11,Address}; end
						4'h7: begin nDat <= 71;  StrtSq <= {2'b11,Address}; end
						4'h8: begin nDat <= 71;  StrtSq <= {2'b11,Address}; end
						4'h9: nDat <= 7;
						4'ha: nDat <= 7;
						4'hb: nDat <= 18;
						4'hc: nDat <= 63;
						4'hd: nDat <= 63;
						4'he: nDat <= 63;
						4'hf: begin nDat <= 7; CalStrobe <= 1'b1; end
					endcase 
				end
		Ct66:	begin
//					$display("%g\t FPGA_DAQ_TKR6:  %b CMDtoChips=%b,  Dout=%b",$time,State,CMDtoChips,Dout);
					Cnt <= Cnt + 1;
					CalStrobe <= 1'b0;
					if (ReadRegCmd && Cnt>0) begin  //This timing to receive register data back may differ between CPU sim vs FPGA board
						case(CmdSav[8:4])			//Select the correct chip from which to receive register data
								5'b00000: StrtSq <= {StrtSq[4:0],Data[0]};         
								5'b00001: StrtSq <= {StrtSq[4:0],Data[1]};
								5'b00010: StrtSq <= {StrtSq[4:0],Data[2]};
								5'b00011: StrtSq <= {StrtSq[4:0],Data[3]};
								5'b00100: StrtSq <= {StrtSq[4:0],Data[4]};
								5'b00101: StrtSq <= {StrtSq[4:0],Data[5]};
						endcase
					end
				end
		RdCm:	begin
					Cnt <= Cnt + 1;
					RegIn <= {RegIn[1:0],CmdIn};		//Shift in the 3-bit local command
				end
		Deco:	begin
					$display("%g\t FPGA_DAQ_TKR6:  local command string=%b",$time,RegIn);
					Parity <= Parity^CmdIn;     	//Including the parity bit in the parity calculation
					Cnt <= 0;
					if (ThisFPGA) begin
						case (RegIn)
							cmdTest: RegOut <= {2'b11,Address,72'b110001011111000001111110000011111100000111111000001111110000011111100011}; 
							cmdStRn: InProg <= 1'b1;
							cmdEnRn: begin
										InProg <= 1'b0;
										EndRun <= 1'b1;
									 end
							cmdRdFg: begin
										RegOut[1:0] <= 2'b11;
										RegOut[17:2] <= NSends;
										RegOut[33:18] <= NReads;
										RegOut[65:34] <= Ntriggers;
										RegOut[77:66] <= {2'b11,Address,4'b1111,TrgErr,Error};      //Start pattern
										Error <= 1'b0;
										$display("%g\t FPGA_DAQ_TKR6: NSends=%d, NReads=%d, Ntriggers=%d",$time,NSends,NReads,Ntriggers);
									 end
							cmdRset: begin
										$display("%g\t FPGA_DAQ_TKR6:  reset command received",$time);
										Reset <= 1'b1;			
									 end
							cmdRsCh: begin
										$display("%g\t FPGA_DAQ_TKR6:  slow reset of ASICs initiated",$time);
										ResetSlow <= 1'b1;		//Reset the ASICs and then reload their configuration
									 end
							cmdSend: begin
//										$display("%g\t FPGA_DAQ_TKR6:  send command received.",$time);
										SendEvt <= 1'b1;		//Trigger the data merger to send out a complete event
										NSends <= NSends + 1;
									 end
						endcase
					end
				end
		WtDn:	begin
					ResetSlow <= 1'b0;			//Long millisecond wait for the reset to complete and amplifiers to settle
				end
		Prty:	begin
					if (Parity) Error <= 1'b1;
					Reset <= 1'b0;
					EndRun <= 1'b0;
					SendEvt <= 1'b0;
				end
		WrWd:	begin
					RegOut <= {RegOut[76:0],1'b0};		//Shifting out the test string or the DAQ counters
					Cnt<=Cnt+1;
				end
	endcase
  end
end

//Matching of the address, either of this chip or the wildcard address
assign ThisFPGA = ((Address==AddrIn || AddrIn==4'hF));

//Recognize when the ASIC command will result in register data coming back
assign ReadRegCmd = (CmdSav[3:0]==4'h3) | (CmdSav[3:0]==4'h4) | (CmdSav[3:0]==4'h5) | (CmdSav[3:0]==4'h6) | (CmdSav[3:0]==4'h7) | (CmdSav[3:0]==4'h8); 

//Program to reset the ASICs without altering their registers
FeReset FeReset_U(DoneRst,CmdRst,Data,ResetSlow,Clock,Reset);

//MUX of the command line going to the chips
always @ (ThisFPGA or CmdIn or State or CmdRst) begin
	if (ThisFPGA && (State == ACmd || State == FeCd || State == Ct66)) CMDtoChips = CmdIn;  //Commands from the event builder
	else if (State == WtDn) CMDtoChips = CmdRst;											//Hand control over to the reset program
	else CMDtoChips = 1'b0;
end

//MUX of the output serial data stream
always @ (State or MuxData or StrtSq or RegOut or ThisFPGA or InProg or ReadRegCmd or Cnt)
begin
	if (InProg) begin
		Dout = MuxData;       												//Event data or TOT calibration data
//	end else if (State == Ct66 && Cnt>0 && ThisFPGA && ReadRegCmd) begin   	//This line for real FPGA
	end else if (State == Ct66 && ThisFPGA && ReadRegCmd) begin    			//This line for cpu sims?
		Dout = StrtSq[5];     												//Register data coming back from the ASICs
	end else if (ThisFPGA && State == WrWd) begin
		Dout = RegOut[77];    												//DAQ counters
	end else begin
		Dout = 1'b0;
	end
end

//Instantiate the DAQ program that merges data from 6 chips
DataMerge6 DataMerge6_U(Clock,Reset,Data,EndRun,UnDoBuf,NoRead,MergeData,Address,SendEvt);

//always @ (posedge Tack) begin
//	$display("%g\t FPGA_DAQ:  Tack signal",$time);
//end

//State machine to insert TOT events into the output stream when the calibration strobe is used
//Some care by the user must be taken not to send a Read command too soon after the strobe, so that this does
//not conflict with the normal event output.
//These TOT events are distinguished from real events by looking at bit 5 of the number of clusters.  That bit
//will be set for these TOT events but never for real events (since 10 is the maximum number of clusters).
//No CRC is attached to the end of these packets.

parameter [7:0] WaitTOT= 8'b00000001; //Wait for a signal that a calibration strobe is starting
parameter [7:0] TReqTOT= 8'b00000010; //Count until the TReq goes high
parameter [7:0] CTOTTOT= 8'b00000100; //Count the TOT, until TReq goes low
parameter [7:0] SOutTOT= 8'b00001000; //Initialize the output sequence, taking over the data output line
parameter [7:0] SHdrTOT= 8'b00010000; //Shift out a 6-bit event header
parameter [7:0] SCluTOT= 8'b00100000; //Shift out 6-bit cluster number, with exactly two "clusters" plus bit 4 set (which isn't used in data taking)
parameter [7:0] STrtTOT= 8'b01000000; //Shift out the 12 bit start counter
parameter [7:0] STOTTOT= 8'b10000000; //Shift out the 12 bit TOT counter.  Zero means that no TReq was encountered.  Release the data output line at the end.
reg [7:0] StateTOT, NextStateTOT;
reg [11:0] CntStrt, CntTOT;
reg [11:0] TOTNclus;
reg [17:0] TOTHeader;
reg [6:0] CntShft;
parameter [11:0] MaxCnt= 12'd255;    //Maximum count allowed

//always @ (posedge Clock) begin
//	$display("%g\t   %b    %b     %b     %d    %d   %d   %b %b %b ",$time,StateTOT,TReqChip,CalStrobe,CntStrt,CntTOT,CntShft,TOTHeader,TOTNclus,MuxData);
//end

always @ (StateTOT or CntStrt or CntTOT or CntShft or TOTHeader or TOTNclus or CalStrobe or TReqChip or MergeData)
begin
	case (StateTOT)
		WaitTOT: 	begin
						MuxData = MergeData;
						if (CalStrobe) NextStateTOT = TReqTOT;
						else NextStateTOT = WaitTOT;
					end
		TReqTOT:	begin
						MuxData = 1'b0;
						if (CntStrt == MaxCnt) NextStateTOT = SOutTOT;  //No TReq found; Send out empty event
						else if (TReqChip) NextStateTOT = CTOTTOT;
						else NextStateTOT = TReqTOT;
					end
		CTOTTOT:	begin
						MuxData = 1'b0;
						if (!TReqChip || CntTOT == MaxCnt) NextStateTOT = SOutTOT;
						else NextStateTOT = CTOTTOT;
					end
		SOutTOT:	begin
						MuxData = 1'b0;
						NextStateTOT = SHdrTOT;
					end
		SHdrTOT:	begin
						if (CntShft == 18) begin
							NextStateTOT = SCluTOT;
							MuxData = TOTNclus[11];
						end else begin
							NextStateTOT = SHdrTOT;
							MuxData = TOTHeader[17];
						end
					end
		SCluTOT:	begin
						if (CntShft == 30) begin
							NextStateTOT = STrtTOT;
							MuxData = CntStrt[11];
						end else begin
							NextStateTOT = SCluTOT;
							MuxData = TOTNclus[11];
						end
					end
		STrtTOT:	begin
						if (CntShft == 42) begin
							NextStateTOT = STOTTOT;
							MuxData = CntTOT[11];
						end else begin
							NextStateTOT = STrtTOT;
							MuxData = CntStrt[11];
						end
					end
		STOTTOT:	begin
						if (CntShft == 54) NextStateTOT = WaitTOT;
						else NextStateTOT = STOTTOT;
						MuxData = CntTOT[11];
					end
		default:	begin
						MuxData = MergeData;
						NextStateTOT = WaitTOT;
					end
	endcase
end

always @ (posedge Clock)
begin
	if (ResetHard) begin
		StateTOT <= WaitTOT;
	end else begin
		StateTOT <= NextStateTOT;
		case (StateTOT)
			WaitTOT: 	begin
							CntStrt <= 0;
							CntTOT <= 0;
						end
			TReqTOT:	begin
							CntStrt <= CntStrt + 1;
						end
			CTOTTOT:	begin
							CntTOT <= CntTOT + 1;
						end
			SOutTOT:	begin
							TOTNclus  <= 12'b010010001111;
							TOTHeader <= {2'b10,Address,12'b111111100001};
							CntShft <= 0;
						end
			SHdrTOT:	begin
							TOTHeader <= {TOTHeader[16:0],1'b0};
							CntShft <= CntShft + 1;
							if (CntShft == 12) TOTNclus <= {TOTNclus[10:0],1'b0};
						end
			SCluTOT:	begin
							TOTNclus <= {TOTNclus[10:0],1'b0};
							CntShft <= CntShft + 1;
							if (CntShft == 18) CntStrt <= {CntStrt[10:0],1'b0};
						end
			STrtTOT:	begin
							CntStrt <= {CntStrt[10:0],1'b0};
							CntShft <= CntShft + 1;
							if (CntShft == 30) CntTOT <= {CntTOT[10:0],1'b0};
						end
			STOTTOT:	begin
							CntTOT <= {CntTOT[10:0],1'b0};
							CntShft <= CntShft + 1;
						end
		endcase
	end
end

endmodule
	